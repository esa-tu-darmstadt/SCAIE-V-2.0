module top(input clk, input rst,

	//AXI instr uncached
	output [31:0] IUC_ARADDR,
	output [1:0] IUC_ARBURST,
	output [3:0] IUC_ARCACHE,
	output [1:0] IUC_ARID,
	output [3:0] IUC_ARLEN,
	output [1:0] IUC_ARLOCK,
	output [2:0] IUC_ARPROT,
	input IUC_ARREADY,
	output [2:0] IUC_ARSIZE,
	output IUC_ARVALID,
	output [31:0] IUC_AWADDR,
	output [1:0] IUC_AWBURST,
	output [3:0] IUC_AWCACHE,
	output [1:0] IUC_AWID,
	output [3:0] IUC_AWLEN,
	output [1:0] IUC_AWLOCK,
	output [2:0] IUC_AWPROT,
	input IUC_AWREADY,
	output [2:0] IUC_AWSIZE,
	output IUC_AWVALID,
	input [1:0] IUC_BID,
	output IUC_BREADY,
	input [1:0] IUC_BRESP,
	input IUC_BVALID,
	input [31:0] IUC_RDATA,
	input [1:0] IUC_RID,
	input IUC_RLAST,
	output IUC_RREADY,
	input [1:0] IUC_RRESP,
	input IUC_RVALID,
	output [31:0] IUC_WDATA,
	output [1:0] IUC_WID,
	output IUC_WLAST,
	input IUC_WREADY,
	output [3:0] IUC_WSTRB,
	output IUC_WVALID,

	//AXI data uncached
	output [31:0] DUC_ARADDR,
	output [1:0] DUC_ARBURST,
	output [3:0] DUC_ARCACHE,
	output [1:0] DUC_ARID,
	output [3:0] DUC_ARLEN,
	output [1:0] DUC_ARLOCK,
	output [2:0] DUC_ARPROT,
	input DUC_ARREADY,
	output [2:0] DUC_ARSIZE,
	output DUC_ARVALID,
	output [31:0] DUC_AWADDR,
	output [1:0] DUC_AWBURST,
	output [3:0] DUC_AWCACHE,
	output [1:0] DUC_AWID,
	output [3:0] DUC_AWLEN,
	output [1:0] DUC_AWLOCK,
	output [2:0] DUC_AWPROT,
	input DUC_AWREADY,
	output [2:0] DUC_AWSIZE,
	output DUC_AWVALID,
	input [1:0] DUC_BID,
	output DUC_BREADY,
	input [1:0] DUC_BRESP,
	input DUC_BVALID,
	input [31:0] DUC_RDATA,
	input [1:0] DUC_RID,
	input DUC_RLAST,
	output DUC_RREADY,
	input [1:0] DUC_RRESP,
	input DUC_RVALID,
	output [31:0] DUC_WDATA,
	output [1:0] DUC_WID,
	output DUC_WLAST,
	input DUC_WREADY,
	output [3:0] DUC_WSTRB,
	output DUC_WVALID,
	
	input global_interrupts,
	input timer_interrupt,
	input [63:0] timer_value);

    //SCAIEV MAKETOP COREWIRES
	
    orca orca_inst(
        .clk(clk), 
        .reset(0), //TODO: Should actually be connected to rst. However, the core converted to a Verilog netlist does not appear to work after reset is asserted..?

		.IUC_ARADDR(IUC_ARADDR),
		.IUC_ARBURST(IUC_ARBURST),
		.IUC_ARCACHE(IUC_ARCACHE),
		.IUC_ARID(IUC_ARID),
		.IUC_ARLEN(IUC_ARLEN),
		.IUC_ARLOCK(IUC_ARLOCK),
		.IUC_ARPROT(IUC_ARPROT),
		.IUC_ARREADY(IUC_ARREADY),
		.IUC_ARSIZE(IUC_ARSIZE),
		.IUC_ARVALID(IUC_ARVALID),
		.IUC_AWADDR(IUC_AWADDR),
		.IUC_AWBURST(IUC_AWBURST),
		.IUC_AWCACHE(IUC_AWCACHE),
		.IUC_AWID(IUC_AWID),
		.IUC_AWLEN(IUC_AWLEN),
		.IUC_AWLOCK(IUC_AWLOCK),
		.IUC_AWPROT(IUC_AWPROT),
		.IUC_AWREADY(IUC_AWREADY),
		.IUC_AWSIZE(IUC_AWSIZE),
		.IUC_AWVALID(IUC_AWVALID),
		.IUC_BID(IUC_BID),
		.IUC_BREADY(IUC_BREADY),
		.IUC_BRESP(IUC_BRESP),
		.IUC_BVALID(IUC_BVALID),
		.IUC_RDATA(IUC_RDATA),
		.IUC_RID(IUC_RID),
		.IUC_RLAST(IUC_RLAST),
		.IUC_RREADY(IUC_RREADY),
		.IUC_RRESP(IUC_RRESP),
		.IUC_RVALID(IUC_RVALID),
		.IUC_WDATA(IUC_WDATA),
		.IUC_WID(IUC_WID),
		.IUC_WLAST(IUC_WLAST),
		.IUC_WREADY(IUC_WREADY),
		.IUC_WSTRB(IUC_WSTRB),
		.IUC_WVALID(IUC_WVALID),

		.DUC_ARADDR(DUC_ARADDR),
		.DUC_ARBURST(DUC_ARBURST),
		.DUC_ARCACHE(DUC_ARCACHE),
		.DUC_ARID(DUC_ARID),
		.DUC_ARLEN(DUC_ARLEN),
		.DUC_ARLOCK(DUC_ARLOCK),
		.DUC_ARPROT(DUC_ARPROT),
		.DUC_ARREADY(DUC_ARREADY),
		.DUC_ARSIZE(DUC_ARSIZE),
		.DUC_ARVALID(DUC_ARVALID),
		.DUC_AWADDR(DUC_AWADDR),
		.DUC_AWBURST(DUC_AWBURST),
		.DUC_AWCACHE(DUC_AWCACHE),
		.DUC_AWID(DUC_AWID),
		.DUC_AWLEN(DUC_AWLEN),
		.DUC_AWLOCK(DUC_AWLOCK),
		.DUC_AWPROT(DUC_AWPROT),
		.DUC_AWREADY(DUC_AWREADY),
		.DUC_AWSIZE(DUC_AWSIZE),
		.DUC_AWVALID(DUC_AWVALID),
		.DUC_BID(DUC_BID),
		.DUC_BREADY(DUC_BREADY),
		.DUC_BRESP(DUC_BRESP),
		.DUC_BVALID(DUC_BVALID),
		.DUC_RDATA(DUC_RDATA),
		.DUC_RID(DUC_RID),
		.DUC_RLAST(DUC_RLAST),
		.DUC_RREADY(DUC_RREADY),
		.DUC_RRESP(DUC_RRESP),
		.DUC_RVALID(DUC_RVALID),
		.DUC_WDATA(DUC_WDATA),
		.DUC_WID(DUC_WID),
		.DUC_WLAST(DUC_WLAST),
		.DUC_WREADY(DUC_WREADY),
		.DUC_WSTRB(DUC_WSTRB),
		.DUC_WVALID(DUC_WVALID),

		.global_interrupts(global_interrupts),
		.timer_interrupt(timer_interrupt),
		.timer_value(timer_value),

		.DC_ARADDR(),
		.DC_ARBURST(),
		.DC_ARCACHE(),
		.DC_ARID(),
		.DC_ARLEN(),
		.DC_ARLOCK(),
		.DC_ARPROT(),
		.DC_ARREADY(),
		.DC_ARSIZE(),
		.DC_ARVALID(),
		.DC_AWADDR(),
		.DC_AWBURST(),
		.DC_AWCACHE(),
		.DC_AWID(),
		.DC_AWLEN(),
		.DC_AWLOCK(),
		.DC_AWPROT(),
		.DC_AWREADY(),
		.DC_AWSIZE(),
		.DC_AWVALID(),
		.DC_BID(),
		.DC_BREADY(),
		.DC_BRESP(),
		.DC_BVALID(),
		.DC_RDATA(),
		.DC_RID(),
		.DC_RLAST(),
		.DC_RREADY(),
		.DC_RRESP(),
		.DC_RVALID(),
		.DC_WDATA(),
		.DC_WID(),
		.DC_WLAST(),
		.DC_WREADY(),
		.DC_WSTRB(),
		.DC_WVALID(),
		.DLMB_AS(),
		.DLMB_Addr(),
		.DLMB_Byte_Enable(),
		.DLMB_CE(),
		.DLMB_Data_Read(),
		.DLMB_Data_Write(),
		.DLMB_Read_Strobe(),
		.DLMB_Ready(),
		.DLMB_UE(),
		.DLMB_Wait(),
		.DLMB_Write_Strobe(),
		.IC_ARADDR(),
		.IC_ARBURST(),
		.IC_ARCACHE(),
		.IC_ARID(),
		.IC_ARLEN(),
		.IC_ARLOCK(),
		.IC_ARPROT(),
		.IC_ARREADY(),
		.IC_ARSIZE(),
		.IC_ARVALID(),
		.IC_AWADDR(),
		.IC_AWBURST(),
		.IC_AWCACHE(),
		.IC_AWID(),
		.IC_AWLEN(),
		.IC_AWLOCK(),
		.IC_AWPROT(),
		.IC_AWREADY(),
		.IC_AWSIZE(),
		.IC_AWVALID(),
		.IC_BID(),
		.IC_BREADY(),
		.IC_BRESP(),
		.IC_BVALID(),
		.IC_RDATA(),
		.IC_RID(),
		.IC_RLAST(),
		.IC_RREADY(),
		.IC_RRESP(),
		.IC_RVALID(),
		.IC_WDATA(),
		.IC_WID(),
		.IC_WLAST(),
		.IC_WREADY(),
		.IC_WSTRB(),
		.IC_WVALID(),
		.ILMB_AS(),
		.ILMB_Addr(),
		.ILMB_Byte_Enable(),
		.ILMB_CE(),
		.ILMB_Data_Read(),
		.ILMB_Data_Write(),
		.ILMB_Read_Strobe(),
		.ILMB_Ready(),
		.ILMB_UE(),
		.ILMB_Wait(),
		.ILMB_Write_Strobe(),
		.avm_data_address(),
		.avm_data_byteenable(),
		.avm_data_read(),
		.avm_data_readdata(),
		.avm_data_readdatavalid(),
		.avm_data_waitrequest(),
		.avm_data_write(),
		.avm_data_writedata(),
		.avm_instruction_address(),
		.avm_instruction_read(),
		.avm_instruction_readdata(),
		.avm_instruction_readdatavalid(),
		.avm_instruction_waitrequest(),
		.data_ACK_I(),
		.data_ADR_O(),
		.data_CTI_O(),
		.data_CYC_O(),
		.data_DAT_I(),
		.data_DAT_O(),
		.data_SEL_O(),
		.data_STALL_I(),
		.data_STB_O(),
		.data_WE_O(),
		.instr_ACK_I(),
		.instr_ADR_O(),
		.instr_CTI_O(),
		.instr_CYC_O(),
		.instr_DAT_I(),
		.instr_STALL_I(),
		.instr_STB_O(),
		.vcp_alu_data1(),
		.vcp_alu_data2(),
		.vcp_alu_result(),
		.vcp_alu_result_valid(),
		.vcp_alu_source_valid(),
		.vcp_data0(),
		.vcp_data1(),
		.vcp_data2(),
		.vcp_illegal(),
		.vcp_instruction(),
		.vcp_ready(),
		.vcp_valid_instr(),
		.vcp_writeback_data(),
		.vcp_writeback_en()

        //SCAIEV MAKETOP COREPINS
    );

    //SCAIEV MAKETOP ISAXWIRES
    
    //SCAIEV MAKETOP SCAL
    
    //SCAIEV MAKETOP ISAXINST
	
endmodule
