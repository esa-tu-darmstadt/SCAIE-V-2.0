module top(input clk, rst,

  input  [3 : 0] set_verbosity_verbosity,
  input  [63 : 0] set_verbosity_logdelay,
  input  EN_set_verbosity,
  output RDY_set_verbosity,

  input  cpu_reset_server_request_put,
  input  EN_cpu_reset_server_request_put,
  output RDY_cpu_reset_server_request_put,

  input  EN_cpu_reset_server_response_get,
  output cpu_reset_server_response_get,
  output RDY_cpu_reset_server_response_get,

  output cpu_imem_master_awvalid,
  output [3 : 0] cpu_imem_master_awid,
  output [63 : 0] cpu_imem_master_awaddr,
  output [7 : 0] cpu_imem_master_awlen,
  output [2 : 0] cpu_imem_master_awsize,
  output [1 : 0] cpu_imem_master_awburst,
  output cpu_imem_master_awlock,
  output [3 : 0] cpu_imem_master_awcache,
  output [2 : 0] cpu_imem_master_awprot,
  output [3 : 0] cpu_imem_master_awqos,
  output [3 : 0] cpu_imem_master_awregion,
  input  cpu_imem_master_awready,
  output cpu_imem_master_wvalid,
  output [63 : 0] cpu_imem_master_wdata,
  output [7 : 0] cpu_imem_master_wstrb,
  output cpu_imem_master_wlast,
  input  cpu_imem_master_wready,
  input  cpu_imem_master_bvalid,
  input  [3 : 0] cpu_imem_master_bid,
  input  [1 : 0] cpu_imem_master_bresp,
  output cpu_imem_master_bready,
  output cpu_imem_master_arvalid,
  output [3 : 0] cpu_imem_master_arid,
  output [63 : 0] cpu_imem_master_araddr,
  output [7 : 0] cpu_imem_master_arlen,
  output [2 : 0] cpu_imem_master_arsize,
  output [1 : 0] cpu_imem_master_arburst,
  output cpu_imem_master_arlock,
  output [3 : 0] cpu_imem_master_arcache,
  output [2 : 0] cpu_imem_master_arprot,
  output [3 : 0] cpu_imem_master_arqos,
  output [3 : 0] cpu_imem_master_arregion,
  input  cpu_imem_master_arready,
  input  cpu_imem_master_rvalid,
  input  [3 : 0] cpu_imem_master_rid,
  input  [63 : 0] cpu_imem_master_rdata,
  input  [1 : 0] cpu_imem_master_rresp,
  input  cpu_imem_master_rlast,
  output cpu_imem_master_rready,

  output cpu_dmem_master_awvalid,
  output [3 : 0] cpu_dmem_master_awid,
  output [63 : 0] cpu_dmem_master_awaddr,
  output [7 : 0] cpu_dmem_master_awlen,
  output [2 : 0] cpu_dmem_master_awsize,
  output [1 : 0] cpu_dmem_master_awburst,
  output cpu_dmem_master_awlock,
  output [3 : 0] cpu_dmem_master_awcache,
  output [2 : 0] cpu_dmem_master_awprot,
  output [3 : 0] cpu_dmem_master_awqos,
  output [3 : 0] cpu_dmem_master_awregion,
  input  cpu_dmem_master_awready,
  output cpu_dmem_master_wvalid,
  output [63 : 0] cpu_dmem_master_wdata,
  output [7 : 0] cpu_dmem_master_wstrb,
  output cpu_dmem_master_wlast,
  input  cpu_dmem_master_wready,
  input  cpu_dmem_master_bvalid,
  input  [3 : 0] cpu_dmem_master_bid,
  input  [1 : 0] cpu_dmem_master_bresp,
  output cpu_dmem_master_bready,
  output cpu_dmem_master_arvalid,
  output [3 : 0] cpu_dmem_master_arid,
  output [63 : 0] cpu_dmem_master_araddr,
  output [7 : 0] cpu_dmem_master_arlen,
  output [2 : 0] cpu_dmem_master_arsize,
  output [1 : 0] cpu_dmem_master_arburst,
  output cpu_dmem_master_arlock,
  output [3 : 0] cpu_dmem_master_arcache,
  output [2 : 0] cpu_dmem_master_arprot,
  output [3 : 0] cpu_dmem_master_arqos,
  output [3 : 0] cpu_dmem_master_arregion,
  input  cpu_dmem_master_arready,
  input  cpu_dmem_master_rvalid,
  input  [3 : 0] cpu_dmem_master_rid,
  input  [63 : 0] cpu_dmem_master_rdata,
  input  [1 : 0] cpu_dmem_master_rresp,
  input  cpu_dmem_master_rlast,
  output cpu_dmem_master_rready,

  input  core_external_interrupt_sources_0_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_1_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_2_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_3_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_4_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_5_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_6_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_7_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_8_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_9_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_10_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_11_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_12_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_13_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_14_m_interrupt_req_set_not_clear,
  input  core_external_interrupt_sources_15_m_interrupt_req_set_not_clear,

  input  nmi_req_set_not_clear);
	
  //SCAIEV MAKETOP COREWIRES
  
    mkCore Piccolo_inst(
        .CLK(clk),
        .RST_N(~rst),

        .set_verbosity_verbosity(set_verbosity_verbosity),
        .set_verbosity_logdelay(set_verbosity_logdelay),
        .EN_set_verbosity(EN_set_verbosity),
        .RDY_set_verbosity(RDY_set_verbosity),

        .cpu_reset_server_request_put(cpu_reset_server_request_put),
        .EN_cpu_reset_server_request_put(EN_cpu_reset_server_request_put),
        .RDY_cpu_reset_server_request_put(RDY_cpu_reset_server_request_put),

        .EN_cpu_reset_server_response_get(EN_cpu_reset_server_response_get),
        .cpu_reset_server_response_get(cpu_reset_server_response_get),
        .RDY_cpu_reset_server_response_get(RDY_cpu_reset_server_response_get),

        .cpu_imem_master_awvalid(cpu_imem_master_awvalid),
        .cpu_imem_master_awid(cpu_imem_master_awid),
        .cpu_imem_master_awaddr(cpu_imem_master_awaddr),
        .cpu_imem_master_awlen(cpu_imem_master_awlen),
        .cpu_imem_master_awsize(cpu_imem_master_awsize),
        .cpu_imem_master_awburst(cpu_imem_master_awburst),
        .cpu_imem_master_awlock(cpu_imem_master_awlock),
        .cpu_imem_master_awcache(cpu_imem_master_awcache),
        .cpu_imem_master_awprot(cpu_imem_master_awprot),
        .cpu_imem_master_awqos(cpu_imem_master_awqos),
        .cpu_imem_master_awregion(cpu_imem_master_awregion),
        .cpu_imem_master_awready(cpu_imem_master_awready),
        .cpu_imem_master_wvalid(cpu_imem_master_wvalid),
        .cpu_imem_master_wdata(cpu_imem_master_wdata),
        .cpu_imem_master_wstrb(cpu_imem_master_wstrb),
        .cpu_imem_master_wlast(cpu_imem_master_wlast),
        .cpu_imem_master_wready(cpu_imem_master_wready),
        .cpu_imem_master_bvalid(cpu_imem_master_bvalid),
        .cpu_imem_master_bid(cpu_imem_master_bid),
        .cpu_imem_master_bresp(cpu_imem_master_bresp),
        .cpu_imem_master_bready(cpu_imem_master_bready),
        .cpu_imem_master_arvalid(cpu_imem_master_arvalid),
        .cpu_imem_master_arid(cpu_imem_master_arid),
        .cpu_imem_master_araddr(cpu_imem_master_araddr),
        .cpu_imem_master_arlen(cpu_imem_master_arlen),
        .cpu_imem_master_arsize(cpu_imem_master_arsize),
        .cpu_imem_master_arburst(cpu_imem_master_arburst),
        .cpu_imem_master_arlock(cpu_imem_master_arlock),
        .cpu_imem_master_arcache(cpu_imem_master_arcache),
        .cpu_imem_master_arprot(cpu_imem_master_arprot),
        .cpu_imem_master_arqos(cpu_imem_master_arqos),
        .cpu_imem_master_arregion(cpu_imem_master_arregion),
        .cpu_imem_master_arready(cpu_imem_master_arready),
        .cpu_imem_master_rvalid(cpu_imem_master_rvalid),
        .cpu_imem_master_rid(cpu_imem_master_rid),
        .cpu_imem_master_rdata(cpu_imem_master_rdata),
        .cpu_imem_master_rresp(cpu_imem_master_rresp),
        .cpu_imem_master_rlast(cpu_imem_master_rlast),
        .cpu_imem_master_rready(cpu_imem_master_rready),

        .cpu_dmem_master_awvalid(cpu_dmem_master_awvalid),
        .cpu_dmem_master_awid(cpu_dmem_master_awid),
        .cpu_dmem_master_awaddr(cpu_dmem_master_awaddr),
        .cpu_dmem_master_awlen(cpu_dmem_master_awlen),
        .cpu_dmem_master_awsize(cpu_dmem_master_awsize),
        .cpu_dmem_master_awburst(cpu_dmem_master_awburst),
        .cpu_dmem_master_awlock(cpu_dmem_master_awlock),
        .cpu_dmem_master_awcache(cpu_dmem_master_awcache),
        .cpu_dmem_master_awprot(cpu_dmem_master_awprot),
        .cpu_dmem_master_awqos(cpu_dmem_master_awqos),
        .cpu_dmem_master_awregion(cpu_dmem_master_awregion),
        .cpu_dmem_master_awready(cpu_dmem_master_awready),
        .cpu_dmem_master_wvalid(cpu_dmem_master_wvalid),
        .cpu_dmem_master_wdata(cpu_dmem_master_wdata),
        .cpu_dmem_master_wstrb(cpu_dmem_master_wstrb),
        .cpu_dmem_master_wlast(cpu_dmem_master_wlast),
        .cpu_dmem_master_wready(cpu_dmem_master_wready),
        .cpu_dmem_master_bvalid(cpu_dmem_master_bvalid),
        .cpu_dmem_master_bid(cpu_dmem_master_bid),
        .cpu_dmem_master_bresp(cpu_dmem_master_bresp),
        .cpu_dmem_master_bready(cpu_dmem_master_bready),
        .cpu_dmem_master_arvalid(cpu_dmem_master_arvalid),
        .cpu_dmem_master_arid(cpu_dmem_master_arid),
        .cpu_dmem_master_araddr(cpu_dmem_master_araddr),
        .cpu_dmem_master_arlen(cpu_dmem_master_arlen),
        .cpu_dmem_master_arsize(cpu_dmem_master_arsize),
        .cpu_dmem_master_arburst(cpu_dmem_master_arburst),
        .cpu_dmem_master_arlock(cpu_dmem_master_arlock),
        .cpu_dmem_master_arcache(cpu_dmem_master_arcache),
        .cpu_dmem_master_arprot(cpu_dmem_master_arprot),
        .cpu_dmem_master_arqos(cpu_dmem_master_arqos),
        .cpu_dmem_master_arregion(cpu_dmem_master_arregion),
        .cpu_dmem_master_arready(cpu_dmem_master_arready),
        .cpu_dmem_master_rvalid(cpu_dmem_master_rvalid),
        .cpu_dmem_master_rid(cpu_dmem_master_rid),
        .cpu_dmem_master_rdata(cpu_dmem_master_rdata),
        .cpu_dmem_master_rresp(cpu_dmem_master_rresp),
        .cpu_dmem_master_rlast(cpu_dmem_master_rlast),
        .cpu_dmem_master_rready(cpu_dmem_master_rready),

        .core_external_interrupt_sources_0_m_interrupt_req_set_not_clear(core_external_interrupt_sources_0_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_1_m_interrupt_req_set_not_clear(core_external_interrupt_sources_1_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_2_m_interrupt_req_set_not_clear(core_external_interrupt_sources_2_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_3_m_interrupt_req_set_not_clear(core_external_interrupt_sources_3_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_4_m_interrupt_req_set_not_clear(core_external_interrupt_sources_4_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_5_m_interrupt_req_set_not_clear(core_external_interrupt_sources_5_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_6_m_interrupt_req_set_not_clear(core_external_interrupt_sources_6_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_7_m_interrupt_req_set_not_clear(core_external_interrupt_sources_7_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_8_m_interrupt_req_set_not_clear(core_external_interrupt_sources_8_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_9_m_interrupt_req_set_not_clear(core_external_interrupt_sources_9_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_10_m_interrupt_req_set_not_clear(core_external_interrupt_sources_10_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_11_m_interrupt_req_set_not_clear(core_external_interrupt_sources_11_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_12_m_interrupt_req_set_not_clear(core_external_interrupt_sources_12_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_13_m_interrupt_req_set_not_clear(core_external_interrupt_sources_13_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_14_m_interrupt_req_set_not_clear(core_external_interrupt_sources_14_m_interrupt_req_set_not_clear),
        .core_external_interrupt_sources_15_m_interrupt_req_set_not_clear(core_external_interrupt_sources_15_m_interrupt_req_set_not_clear),

        .nmi_req_set_not_clear(nmi_req_set_not_clear)

        //SCAIEV MAKETOP COREPINS
    );

    //SCAIEV MAKETOP ISAXWIRES
    
    //SCAIEV MAKETOP SCAL
    
    //SCAIEV MAKETOP ISAXINST
	
endmodule
