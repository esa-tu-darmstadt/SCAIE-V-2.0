module cva5_top (
    input wire clk,
    input wire rst,

	output wire [31:0] instruction_bram_addr,
	output wire        instruction_bram_en,
	output wire [3:0]  instruction_bram_we,
	output wire [31:0] instruction_bram_din,
	input  wire [31:0] instruction_bram_dout,

	output wire [31:0] data_bram_addr,
	output wire        data_bram_en,
	output wire [3:0]  data_bram_we,
	output wire [31:0] data_bram_din,
	input  wire [31:0] data_bram_dout,
    
    // Generic LSU memory interface
    output wire dgeneric_new_request,
    output wire [31:0] dgeneric_addr,
    output wire dgeneric_re,
    output wire dgeneric_we,
    output wire [3:0] dgeneric_be,
    output wire [31:0] dgeneric_data_in,
    input wire [31:0] dgeneric_data_out,
    input wire dgeneric_data_valid,
    input wire dgeneric_ready,

    // Generic Fetch memory interface
    output wire igeneric_new_request,
    output wire [31:0] igeneric_addr,
    output wire igeneric_re,
    output wire igeneric_we,
    output wire [3:0] igeneric_be,
    output wire [31:0] igeneric_data_in,
    input wire [31:0] igeneric_data_out,
    input wire igeneric_data_valid,
    input wire igeneric_ready,

	// AXI Bus
	// AXI Write Channels
	output wire                            m_axi_awvalid,
	input  wire                            m_axi_awready,
	output wire [5:0]                      m_axi_awid,
	output wire [31:0]                     m_axi_awaddr,
	//~ output wire [3:0]                      m_axi_awregion,
	output wire [7:0]                      m_axi_awlen,
	output wire [2:0]                      m_axi_awsize,
	output wire [1:0]                      m_axi_awburst,
	//~ output wire                            m_axi_awlock,
	output wire [3:0]                      m_axi_awcache,
	//~ output wire [2:0]                      m_axi_awprot,
	//~ output wire [3:0]                      m_axi_awqos,

	output wire                            m_axi_wvalid,
	input  wire                            m_axi_wready,
	output wire [31:0]                     m_axi_wdata,
	output wire [3:0]                      m_axi_wstrb,
	output wire                            m_axi_wlast,

	input  wire                            m_axi_bvalid,
	output wire                            m_axi_bready,
	input  wire [1:0]                      m_axi_bresp,
	input  wire [5:0]                      m_axi_bid,

	// AXI Read Channels
	output wire                            m_axi_arvalid,
	input  wire                            m_axi_arready,
	output wire [5:0]                      m_axi_arid,
	output wire [31:0]                     m_axi_araddr,
	//~ output wire [3:0]                      m_axi_arregion,
	output wire [7:0]                      m_axi_arlen,
	output wire [2:0]                      m_axi_arsize,
	output wire [1:0]                      m_axi_arburst,
	//~ output wire                            m_axi_arlock,
	output wire [3:0]                      m_axi_arcache,
	//~ output wire [2:0]                      m_axi_arprot,
	//~ output wire [3:0]                      m_axi_arqos,

	input  wire                            m_axi_rvalid,
	output wire                            m_axi_rready,
	input  wire [5:0]                      m_axi_rid,
	input  wire [31:0]                     m_axi_rdata,
	input  wire [1:0]                      m_axi_rresp,
	input  wire                            m_axi_rlast,

	// AXI Cache
	// AXI Write Channels
	output wire                            m_axi_cache_awvalid,
	input  wire                            m_axi_cache_awready,
	output wire [5:0]                      m_axi_cache_awid,
	output wire [31:0]                     m_axi_cache_awaddr,
	//~ output wire [3:0]                      m_axi_cache_awregion,
	output wire [7:0]                      m_axi_cache_awlen,
	output wire [2:0]                      m_axi_cache_awsize,
	output wire [1:0]                      m_axi_cache_awburst,
	//~ output wire                            m_axi_cache_awlock,
	output wire [3:0]                      m_axi_cache_awcache,
	output wire [2:0]                      m_axi_cache_awprot,
	//~ output wire [3:0]                      m_axi_cache_awqos,

	output wire                            m_axi_cache_wvalid,
	input  wire                            m_axi_cache_wready,
	output wire [31:0]                     m_axi_cache_wdata,
	output wire [3:0]                      m_axi_cache_wstrb,
	output wire                            m_axi_cache_wlast,

	input  wire                            m_axi_cache_bvalid,
	output wire                            m_axi_cache_bready,
	input  wire [1:0]                      m_axi_cache_bresp,
	input  wire [5:0]                      m_axi_cache_bid,

	// AXI Read Channels
	output wire                            m_axi_cache_arvalid,
	input  wire                            m_axi_cache_arready,
	output wire [5:0]                      m_axi_cache_arid,
	output wire [31:0]                     m_axi_cache_araddr,
	//~ output wire [3:0]                      m_axi_cache_arregion,
	output wire [7:0]                      m_axi_cache_arlen,
	output wire [2:0]                      m_axi_cache_arsize,
	output wire [1:0]                      m_axi_cache_arburst,
	//~ output wire                            m_axi_cache_arlock,
	output wire [3:0]                      m_axi_cache_arcache,
	output wire [2:0]                      m_axi_cache_arprot,
	//~ output wire [3:0]                      m_axi_cache_arqos,

	input  wire                            m_axi_cache_rvalid,
	output wire                            m_axi_cache_rready,
	input  wire [5:0]                      m_axi_cache_rid,
	input  wire [31:0]                     m_axi_cache_rdata,
	input  wire [1:0]                      m_axi_cache_rresp,
	input  wire                            m_axi_cache_rlast,
	
	input wire timer_interrupt,
	input wire interrupt
);

    //SCAIEV MAKETOP COREWIRES

	assign dgeneric_new_request = 0;
	assign igeneric_new_request = 0;
    cva5_wrapper cva5 (
        .clk(clk),
        .rst(rst),

        .instruction_bram_addr(instruction_bram_addr),
        .instruction_bram_en(instruction_bram_en),
        .instruction_bram_we(instruction_bram_we),
        .instruction_bram_din(instruction_bram_din),
        .instruction_bram_dout(instruction_bram_dout),
        .data_bram_addr(data_bram_addr),
        .data_bram_en(data_bram_en),
        .data_bram_we(data_bram_we),
        .data_bram_din(data_bram_din),
        .data_bram_dout(data_bram_dout),
        .m_axi_awvalid(m_axi_awvalid),
        .m_axi_awready(m_axi_awready),
        .m_axi_awid(m_axi_awid),
        .m_axi_awaddr(m_axi_awaddr),
        //.m_axi_awregion(m_axi_awregion),
        .m_axi_awlen(m_axi_awlen),
        .m_axi_awsize(m_axi_awsize),
        .m_axi_awburst(m_axi_awburst),
        //.m_axi_awlock(m_axi_awlock),
        .m_axi_awcache(m_axi_awcache),
        //.m_axi_awprot(m_axi_awprot),
        //.m_axi_awqos(m_axi_awqos),
        .m_axi_wvalid(m_axi_wvalid),
        .m_axi_wready(m_axi_wready),
        .m_axi_wdata(m_axi_wdata),
        .m_axi_wstrb(m_axi_wstrb),
        .m_axi_wlast(m_axi_wlast),
        .m_axi_bvalid(m_axi_bvalid),
        .m_axi_bready(m_axi_bready),
        .m_axi_bresp(m_axi_bresp),
        .m_axi_bid(m_axi_bid),
        .m_axi_arvalid(m_axi_arvalid),
        .m_axi_arready(m_axi_arready),
        .m_axi_arid(m_axi_arid),
        .m_axi_araddr(m_axi_araddr),
        //.m_axi_arregion(m_axi_arregion),
        .m_axi_arlen(m_axi_arlen),
        .m_axi_arsize(m_axi_arsize),
        .m_axi_arburst(m_axi_arburst),
        //.m_axi_arlock(m_axi_arlock),
        .m_axi_arcache(m_axi_arcache),
        //.m_axi_arprot(m_axi_arprot),
        //.m_axi_arqos(m_axi_arqos),
        .m_axi_rvalid(m_axi_rvalid),
        .m_axi_rready(m_axi_rready),
        .m_axi_rid(m_axi_rid),
        .m_axi_rdata(m_axi_rdata),
        .m_axi_rresp(m_axi_rresp),
        .m_axi_rlast(m_axi_rlast),

        .axi_awvalid(m_axi_cache_awvalid),
        .axi_awready(m_axi_cache_awready),
        .axi_awid(m_axi_cache_awid),
        .axi_awaddr(m_axi_cache_awaddr),
        .axi_awlen(m_axi_cache_awlen),
        .axi_awsize(m_axi_cache_awsize),
        .axi_awburst(m_axi_cache_awburst),
        .axi_awcache(m_axi_cache_awcache),
        .axi_awprot(m_axi_cache_awprot),
        .axi_wvalid(m_axi_cache_wvalid),
        .axi_wready(m_axi_cache_wready),
        .axi_wdata(m_axi_cache_wdata),
        .axi_wstrb(m_axi_cache_wstrb),
        .axi_wlast(m_axi_cache_wlast),
        .axi_bvalid(m_axi_cache_bvalid),
        .axi_bready(m_axi_cache_bready),
        .axi_bresp(m_axi_cache_bresp),
        .axi_bid(m_axi_cache_bid),
        .axi_arvalid(m_axi_cache_arvalid),
        .axi_arready(m_axi_cache_arready),
        .axi_arid(m_axi_cache_arid),
        .axi_araddr(m_axi_cache_araddr),
        .axi_arlen(m_axi_cache_arlen),
        .axi_arsize(m_axi_cache_arsize),
        .axi_arburst(m_axi_cache_arburst),
        .axi_arcache(m_axi_cache_arcache),
        .axi_arprot(m_axi_cache_arprot),
        .axi_rvalid(m_axi_cache_rvalid),
        .axi_rready(m_axi_cache_rready),
        .axi_rid(m_axi_cache_rid),
        .axi_rdata(m_axi_cache_rdata),
        .axi_rresp(m_axi_cache_rresp),
        .axi_rlast(m_axi_cache_rlast),

        .timer_interrupt(timer_interrupt),
        .interrupt(interrupt)
        
        //SCAIEV MAKETOP COREPINS
    );

    //SCAIEV MAKETOP ISAXWIRES
    
    //SCAIEV MAKETOP SCAL
    
    //SCAIEV MAKETOP ISAXINST

endmodule
